module process

pub const err_not_found = error('The port is available:')

pub const err_command_not_found = error('The executable is not found:')
