module process

pub fn find_process_by_port(port int) ?&Process {
	println(port)
}
