module process

struct Process {
pub:
	proto string
	addr  string
	pid   int
}
