module process

pub fn kill(pid int) ? {
}
